class sequence_item extends uvm_sequence_item;
     `uvm_object_utils(sequence_item)

rand bit rst_n, load;
rand bit [7:0] data_i ; 


logic serial_o ;



endclass //sequence_item extends superClass