package yapp_pkg;

   import uvm_pkg::*;
`include "uvm_macros.svh"

`include "../sv/yapp_packet.sv" 
endpackage




