//`timescale 1ns/1ns

class mem_driver extends uvm_driver#(mem_sequencer_item);
     `uvm_component_utils(mem_driver)

 virtual mem_intf vif ; 
 mem_sequencer_item item ; 
 
 //--------------------------------------------------------
  //Constructor
  //--------------------------------------------------------
  function new(string name = "mem_driver", uvm_component parent);
    super.new(name, parent);
    `uvm_info("DRIVER_CLASS", "Inside Constructor!", UVM_HIGH)
  endfunction: new
  
  
  //--------------------------------------------------------
  //Build Phase
  //--------------------------------------------------------
  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    `uvm_info("DRIVER_CLASS", "Build Phase!", UVM_HIGH)
    
    if(!(uvm_config_db #(virtual mem_intf)::get(this, "*", "vif", vif))) begin
      `uvm_error("DRIVER_CLASS", "Failed to get VIF from config DB!")
    end
    
  endfunction: build_phase
  
  
  //--------------------------------------------------------
  //Connect Phase
  //--------------------------------------------------------
  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    `uvm_info("DRIVER_CLASS", "Connect Phase!", UVM_HIGH)
    
  endfunction: connect_phase
  
  
  //--------------------------------------------------------
  //Run Phase
  //--------------------------------------------------------
  task run_phase (uvm_phase phase);
    super.run_phase(phase);
    `uvm_info("DRIVER_CLASS", "Inside Run Phase!", UVM_HIGH)
    clear();


    forever begin
      @(negedge vif.clk);
      item = mem_sequencer_item::type_id::create("item"); 
      seq_item_port.get_next_item(item);
         `uvm_info("DRIVER_CLASS", "Got transaction from the sequencer!", UVM_LOW)
        vif.addr <= item.addr;
        vif.data_in <= item.data_in;
        vif.read <= item.read;
        vif.write <= item.write;


      seq_item_port.item_done();
    end
    
  endtask: run_phase
  
  
task  clear();
  for (int i =0 ;i<32 ;i++ ) begin
      vif.addr <=i;
        vif.data_in <= 0;
        vif.read <= 0;
        vif.write <= 1;
  end


endtask //


endclass //mem_driver extends superClass