interface piso_intf(input  logic clk);
    
logic rst_n,load;
logic [7:0] data_i; 
logic serial_o;


endinterface //piso_intf