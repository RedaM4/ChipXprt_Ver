interface dut_if(input clk);
    
    logic [7:0] a,b,sum;
    logic carry  ; 

endinterface //dut_if