interface dut_if(input clk);
    logic reset,cmd;
    logic[7:0] addr,data ; 


endinterface //dut_if